
 This is a dummy sv file.

